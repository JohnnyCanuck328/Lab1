library verilog;
use verilog.vl_types.all;
entity eightBitLeftShift_vlg_vec_tst is
end eightBitLeftShift_vlg_vec_tst;
