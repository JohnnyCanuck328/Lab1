library verilog;
use verilog.vl_types.all;
entity controlLogic_vlg_vec_tst is
end controlLogic_vlg_vec_tst;
