library verilog;
use verilog.vl_types.all;
entity eightBitAdder_vlg_vec_tst is
end eightBitAdder_vlg_vec_tst;
