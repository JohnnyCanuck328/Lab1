library verilog;
use verilog.vl_types.all;
entity lab1_vlg_check_tst is
    port(
        NOToutput0      : in     vl_logic;
        NOToutput1      : in     vl_logic;
        NOToutput2      : in     vl_logic;
        NOToutput3      : in     vl_logic;
        NOToutput4      : in     vl_logic;
        NOToutput5      : in     vl_logic;
        NOToutput6      : in     vl_logic;
        NOToutput7      : in     vl_logic;
        output0         : in     vl_logic;
        output1         : in     vl_logic;
        output2         : in     vl_logic;
        output3         : in     vl_logic;
        output4         : in     vl_logic;
        output5         : in     vl_logic;
        output6         : in     vl_logic;
        output7         : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end lab1_vlg_check_tst;
