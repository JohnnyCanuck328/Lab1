library verilog;
use verilog.vl_types.all;
entity dFF_2_vlg_check_tst is
    port(
        o_q             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end dFF_2_vlg_check_tst;
