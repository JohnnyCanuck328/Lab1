library verilog;
use verilog.vl_types.all;
entity h2InMux_vlg_vec_tst is
end h2InMux_vlg_vec_tst;
