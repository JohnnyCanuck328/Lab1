library verilog;
use verilog.vl_types.all;
entity enARdFF_2_vlg_vec_tst is
end enARdFF_2_vlg_vec_tst;
