library verilog;
use verilog.vl_types.all;
entity fourMux_vlg_vec_tst is
end fourMux_vlg_vec_tst;
