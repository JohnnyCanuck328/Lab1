library verilog;
use verilog.vl_types.all;
entity eightbitshiftregister_vlg_vec_tst is
end eightbitshiftregister_vlg_vec_tst;
