library verilog;
use verilog.vl_types.all;
entity dFF_2_vlg_vec_tst is
end dFF_2_vlg_vec_tst;
